module multipliermod(a, b, out);

input [4:0] a;

input [4:0] b;

output [9:0] out;

assign out=(a*b);

endmodule
